`define formatSFP 9
`define exponent 4
`define significand 4


`define SFPWIDTH `formatSFP
`define EXPWIDTH `exponent
`define SIGWIDTH `significand
`define LOW_EXPAND 2
`define FIXWIDTH 21